module _inv(a,y);
input a;		//one input
output y;	//one output

assign y=~a;// y = NOT a	
endmodule	//end of module
